package FIFO_shared_pkg;
	// signal  will assert at the end of the test
	logic test_finished = 0;

	// Define correct and error counters 
	integer correct_count = 0;
	integer error_count = 0;
endpackage 


